module synapse_connection 
#(
	NUM_AXONS = 256,
	NUM_NEURONS = 256
)
(
	input clk,
	input rst,
	input [$clog2(NUM_AXONS)-1:0] axon_number,
    input enable,
	
	output reg synap_con_done,
	output reg [$clog2(NUM_NEURONS)-1:0] neuron_number,
	output reg neuron_number_valid // if that neuron has a connection with the axon spike

);
    wire matrix_connection;
    reg [$clog2(NUM_NEURONS)-1:0] counter;
    
    synap_matrix 
	#(
		.NUM_AXONS(NUM_AXONS),
		.NUM_NEURONS(NUM_AXONS)
	) synap_matrix 
    (
        .clk(clk),
        .rst(rst),
        .axon_number(axon_number),
        .neuron_number(counter),

        .matrix_connection(matrix_connection)
    );

    // // output logic
    // always @(posedge clk) begin
    //     if (rst) begin
    //         neuron_number <= 1'b0;
    //         neuron_number_valid <= 1'b0;
    //     end
    //     else if (enable) begin
    //         if (matrix_connection) begin
    //             neuron_number <= counter;
    //             neuron_number_valid <= 1'b1;
    //         end
    //         else begin 
    //             neuron_number <= 1'b0;
    //             neuron_number_valid <= 1'b0;
    //         end
    //     end
    //     else begin 
    //         neuron_number <= 1'b0;
    //         neuron_number_valid <= 1'b0;
    //     end
    // end

    // // neuron number counter
    // always @(posedge clk) begin
    //     if (rst) begin
    //         counter <= 'b0;
	// 		synap_con_done <= 1'b0;
    //     end
    //     else if (enable) begin 
    //         if (counter == 255) begin
    //             counter <= 1'b0;
    //             synap_con_done <= 1'b1;
    //         end
    //         else begin
    //             counter <= counter + 1'b1;
    //             synap_con_done <= 1'b0;
    //         end
    //     end 
    //     else begin
    //         counter <= counter;
    //         synap_con_done <= 1'b0;
    //     end
    // end

    // counter logic
    always @(posedge clk) begin
        if (rst) begin
            counter <= {($clog2(NUM_AXONS)+1){1'b1}};
        end
        else if (enable) begin
            if (!connection) begin 
                counter <= counter + 1'b1;
            end
            else begin
                counter <= counter;
            end
        end
        else if (synap_con_done) begin
            counter <= {($clog2(NUM_AXONS)+1){1'b1}};
        end
        else begin
            counter <= counter;
        end
    end

    // connection 
    wire connection;
    assign connection = neuron_number_valid ? 1'b0 : matrix_connection;

    // connection & neuron num logic
    always @(posedge clk) begin
        if (rst) begin
            neuron_number <= 1'b0;
            neuron_number_valid <= 1'b0;            
        end
        else if (matrix_connection) begin
            neuron_number <= counter;
            neuron_number_valid <= 1'b1;
        end
        else begin 
            neuron_number <= 1'b0;
            neuron_number_valid <= 1'b0;
        end
    end
    
    // done logic
    always @(posedge clk) begin
        if (rst) begin
			synap_con_done <= 1'b0;
        end
        else if (counter == 256) begin
            synap_con_done <= 1'b1;
        end
        else begin
            synap_con_done <= 1'b0;
        end
    end
    
endmodule

module synap_matrix
#(
	parameter NUM_AXONS = 256,
	parameter NUM_NEURONS = 256,
    parameter bit [0:NUM_NEURONS-1][0:3][63:0] LUT_INIT  = 
    {
        {
        64'hba502b6aaaac7467,
        64'hda869ec794438a23,
        64'h34da925752a6d292,
        64'heaafeaaa292b002b
        },
        {
        64'h8aab130a2029a5b7,
        64'h990ea12ea9afaaae,
        64'hd05bd14ba94b890a,
        64'h9aba2aa960a3aaaa
        },
        {
        64'ha9542152e952658b,
        64'h5893da96bad7a356,
        64'hd65d52585056d032,
        64'heaac24a955a7540c
        },
        {
        64'ha952bd53a8ee4e99,
        64'ha5aa2de8aadbaad6,
        64'h116ca42d86ada32f,
        64'h0aae6ed23df59d62
        },
        {
        64'h928653092aa86695,
        64'h8683a6a2b687b6b3,
        64'h34908497a0cba6c7,
        64'h2aa2e8a840aa50a2
        },
        {
        64'h551bd529b0afbfee,
        64'ha2772ade6ac3e84a,
        64'h50acc2aa82ab10aa,
        64'h6aa91245d4035203
        },
        {
        64'h82a810a1d7773a6c,
        64'hbe4baa6baa2b60aa,
        64'h904ac04af65b325b,
        64'haa8d2aa9a4a9904a
        },
        {
        64'hac502aa96aaa720b,
        64'ha8a828a926983451,
        64'h2a0baa4b2143712b,
        64'h5c462b24aa76ea63
        },
        {
        64'hca1b682b2eaff1c2,
        64'ha90e2446a6db2683,
        64'h206ba46ba82bab2b,
        64'h4aace22aa92f28ee
        },
        {
        64'ha0a82aab2aa926fa,
        64'h95a7b4aea883a54a,
        64'h4aa2ab4ab74ab56f,
        64'h055d91549a538bba
        },
        {
        64'ha128ac2aaaae945e,
        64'hc292828a9232048a,
        64'ha8cb869292839a82,
        64'hcaa32aaa2b4ba14a
        },
        {
        64'ha953215aaa2344ea,
        64'h2db7a5aba8afa27e,
        64'h546bd24baa0b092b,
        64'haaab6aab7502f517
        },
        {
        64'ha952ab50a94257ba,
        64'h5ebab296b696bb52,
        64'h568a504b5157d89f,
        64'heaafa5abd4b6d4be
        },
        {
        64'h20572ab7aaaa5665,
        64'h2aaaa2acb4142156,
        64'h24adb0adba48a94b,
        64'heaab6a5629d422a4
        },
        {
        64'h9483d28b2aa8dae8,
        64'ha00bb04a942394a2,
        64'h28afa957a9172917,
        64'h8aaa824a304b80ab
        },
        {
        64'h122b5e69aea98e5f,
        64'haa4bcb4adb0bc3ab,
        64'h2c11a4aeb8ababae,
        64'heaaaeac8a9cead47
        },
        {
        64'hb4ba968a17d02a3f,
        64'h9a7baa3aa9ba28ba,
        64'ha78aa47bb07b3cfb,
        64'haaa26aaba829a84a
        },
        {
        64'ha851aaa8aaabff90,
        64'ha1a8a56d29d5b151,
        64'h282b8cab86afa4a9,
        64'h90006e17a956aa57
        },
        {
        64'h855a69da2aa802ee,
        64'h9b465246db035142,
        64'h1082a0aba22b3b4b,
        64'h2aacebab3d423553
        },
        {
        64'haa4baa2baaa9a0d5,
        64'h92b390b2a5922a42,
        64'h84968602a61712b7,
        64'h12bd76ab802b84db
        },
        {
        64'ha9412a682aac0cf5,
        64'h925295528512d392,
        64'h0b0f88aa828a92c3,
        64'h2aacaaa8ab522953
        },
        {
        64'ha82b2c28a1288373,
        64'h1a2f092aa923292e,
        64'h602bf32ba9aaaa8a,
        64'h7aa12aa86cabe42b
        },
        {
        64'h2d5535516d4017cd,
        64'h54b6a8928b57a315,
        64'h56d75654569656b7,
        64'hcaad6daa95ae548c
        },
        {
        64'hab46aad3aaab22ef,
        64'haf22a4aea10fa562,
        64'h34a5b4ac92a80b4a,
        64'h8aa924122d45a4b5
        },
        {
        64'h8a8a8aa922aa7c8c,
        64'h95c2b0ca828cd28b,
        64'h08aaa8aba82ab55a,
        64'heaaf6a8305a30a9a
        },
        {
        64'h4aab8aa92aa4ea83,
        64'haa8ac102d52bd2ab,
        64'ha953a853a803aa93,
        64'h8aa8a8a92aabac8a
        },
        {
        64'h8aad9a8d56962c66,
        64'h5257c9d699569b42,
        64'h282b900ad1520352,
        64'h6aa06aab2f2b0b2a
        },
        {
        64'ha8952aab6aae3e74,
        64'hacaca9e52db5b195,
        64'h2b4ba92b810a2ca8,
        64'h7414ac04aab62a4a
        },
        {
        64'hfc6a6a69aaae1696,
        64'hd05652569ad275de,
        64'h161b920bba4bb243,
        64'haaafe82a952a262a
        },
        {
        64'ha54a2aabaaae009f,
        64'h892ba1a2a9aba572,
        64'hc09b83d3a5523147,
        64'he15f105382d70893
        },
        {
        64'hb82bb7a92a270cab,
        64'hb66abe6aadaa20aa,
        64'h280fa8cea4cbb643,
        64'h82a82aaa8a53a822
        },
        {
        64'hb253b14ba3289be3,
        64'h390ee9aea91f2097,
        64'h546bd26b2a6ba909,
        64'h2aa12babf12395ae
        },
        {
        64'ha1aaa02be8a513a3,
        64'h206ba12a812b2126,
        64'he91549456d6a696a,
        64'haaa56aa28b568b57
        },
        {
        64'habd22d532d6f46fb,
        64'hadcaa502a597a196,
        64'h932c83ac81ac392a,
        64'hcaaa6356b724b568
        },
        {
        64'hca5b4229ebafecf0,
        64'hd557ac07aa12aa93,
        64'h3960b56b951b1419,
        64'hcaad4aa9b2aab2ab
        },
        {
        64'h49da49282ead9cdd,
        64'hab5ae9626d26cd92,
        64'hd4e3d4ba968aaa4e,
        64'h0aab0faec76f744a
        },
        {
        64'hc555955755562e7c,
        64'h892388abaaabaaab,
        64'h3153d552c0828803,
        64'h2aa1eaaaaaaabd4b
        },
        {
        64'haa55baab2aab84e4,
        64'haaa928a92d552950,
        64'h282aa92a88938888,
        64'hf450bd4a2a0ae86a
        },
        {
        64'he92b29aaaaa9d89e,
        64'hd52a436a826b666a,
        64'h229a98d3e2d3b92a,
        64'h8aadaaabab7a22db
        },
        {
        64'ha5a82aab2aaabc9b,
        64'hb1578906a8a3a5a2,
        64'h14abaa93a8d73556,
        64'h564bd45ad69750b7
        },
        {
        64'ha929b42baaaca8f0,
        64'hb28b32cab60ba46a,
        64'h288aa28a26cbb28a,
        64'haaacaaaaa84ba84a
        },
        {
        64'hb2a895aaa1aac80e,
        64'h9bafa9aeadaea3af,
        64'hc24bf26bba7a8bb9,
        64'hdaa22aa96a632a0a
        },
        {
        64'hb253aa512942cf8b,
        64'h5abbd4b69497b495,
        64'hd24a5b5b5b52cb16,
        64'h4aafaea0549752e4
        },
        {
        64'h94aaaa8da96ff8f3,
        64'ha92a892c8d2f95b4,
        64'hb697a0b4932ca12a,
        64'h4aaee1592a45b055
        },
        {
        64'h9a6e52a8aaacb0b8,
        64'h99dabeea9e6bd26b,
        64'h2b2ab303bb6a9b9b,
        64'h2aaecaabeb4a8a4a
        },
        {
        64'h50eaeee922ab8cb1,
        64'haa5eea564acad54b,
        64'h20a6b2afbaab224b,
        64'heaa895cc145a1853
        },
        {
        64'hea96155755542430,
        64'hc90a892aaa2a2aab,
        64'h2b4bc552d153c882,
        64'h2aab2aaa24aa354a
        },
        {
        64'haab12aa96aaf10e3,
        64'h9084a04131509a91,
        64'ha9aaa1aab4b3928d,
        64'h9d15b9ec29a629aa
        },
        {
        64'hac72817aaaa83fba,
        64'hb953514e94aa54ab,
        64'h0a4b8b4b895b496a,
        64'h4aaaab999c1b1242
        },
        {
        64'hab4a2b2a6aa1bbea,
        64'h9546950a9aab8a6a,
        64'ha173a157a5571542,
        64'h46aa30ab8aaa8a0b
        },
        {
        64'ha9aa27a82a2a62bf,
        64'hb67a3e6abc2b30ab,
        64'h2a5aa8be34fbb6da,
        64'h0aae2aaa2a3b2ab3
        },
        {
        64'hadab2ca8212e2493,
        64'h9bae89aaa98228aa,
        64'h564ad22abaab8ba8,
        64'haa9eeaa8ee4baa0a
        },
        {
        64'ha428b14868cbdfb2,
        64'h424ab2aa92aaf0ab,
        64'haaa440b55517d556,
        64'h8aa9aaab3aaaf2ac
        },
        {
        64'h245baac72aaff45d,
        64'ha82eb4a4a485200b,
        64'h24a4a4a8a8292a4b,
        64'h6aadaa5728542815
        },
        {
        64'h90974aaa2aa952c4,
        64'hfcd2a8c8a821d286,
        64'ha8a8a8ab815a1946,
        64'h6aacca80114a10ea
        },
        {
        64'h158b95ab3eae738a,
        64'hda56da4a522ad602,
        64'h92d2929782969057,
        64'h2aa818cca8d63053
        },
        {
        64'ha92929674d52dc42,
        64'h90da90dbaa6baa4a,
        64'h4242c3dbc6029183,
        64'h8aa52aabaaaa242b
        },
        {
        64'habd9aaa82aa8cdbf,
        64'h94b4a9953595ac55,
        64'h2a5b9d6f9496d6b4,
        64'hb036a5a528aaba56
        },
        {
        64'h906e962aaeaa3a9c,
        64'hd00b465a921e43f7,
        64'h9ad38adb8a43e92b,
        64'h0aac686b29470a93
        },
        {
        64'ha26b2aa8aaa9fee9,
        64'hb457b4d6accba4ea,
        64'h68aba89aa84ea416,
        64'hc7da34b790aa3aae
        },
        {
        64'h8249822aeaab0caf,
        64'hda828aea92279c02,
        64'h8a5792b612b78ab6,
        64'h4aa9eaa9211aa812
        },
        {
        64'h124a9b1a212c40fc,
        64'haab6aa9ea64bb24e,
        64'h859ba18baaaaabab,
        64'h7abeeaa120b36496
        },
        {
        64'haaa36ad0a94671ae,
        64'h4d2aa982ab036aa8,
        64'hd0ec55945105d943,
        64'h8aa56aa82aa9caae
        },
        {
        64'ha1d72e13a928c0b2,
        64'h292bab2295219530,
        64'h1142886d812d092f,
        64'h0aad6b52a045214c
        },
        {
        64'h88115b08aaaf2091,
        64'hac57a852aa538a53,
        64'hb429966ad53bf54b,
        64'heaa90caab5abb4ab
        },
        {
        64'h148a94ba3ea89484,
        64'hd2d6d29252d3564a,
        64'h20d5a577803714d3,
        64'h6aa0d65acad70257
        },
        {
        64'hc6ab96a99752c032,
        64'haa6bab2aa8aa90ba,
        64'h280aaccaaa4a2a4a,
        64'he29d6aa9a808a8ca
        },
        {
        64'h2ad5aaaa2aaded85,
        64'h8494949113cd3745,
        64'h2aaaa86ab95e1894,
        64'hd1527541212b3aab
        },
        {
        64'hb542e5192eab4d84,
        64'h90a760828053155a,
        64'h14538252aa2bbbab,
        64'hcaa9aaa9254b9552
        },
        {
        64'h294a2a2a6aaf50da,
        64'h91769536acd2ab4a,
        64'h42aec2aab2aeb2a7,
        64'h44bad791166f88af
        },
        {
        64'h8541094baaad81c2,
        64'hc222852a812badc3,
        64'h015684578297d2ab,
        64'hcaa9aaaa3b2228d3
        },
        {
        64'h296b2b4aa92c4f35,
        64'h321b9a7aab63ab2b,
        64'h152bb12baaaaaa8b,
        64'h8ab7ea28bdab702a
        },
        {
        64'hac2d6852e8cea1f2,
        64'h420ba2aaa2aae228,
        64'h98b254965557c046,
        64'haaa5aaa9aaab4ab2
        },
        {
        64'haa55a554a8ec04b7,
        64'hb6533495b49724d4,
        64'h093aacaf94a41497,
        64'h4aaab546b561bc68
        },
        {
        64'h82e7d29aaaade4b2,
        64'ha7d7aed7a2808a83,
        64'haa2aaa2ba9521512,
        64'h8aad62a0961a0e2a
        },
        {
        64'h53fabaa82eafedd5,
        64'ha946eb525a52d34a,
        64'h832b8b23892bab42,
        64'h0aaec769cd0b9323
        },
        {
        64'hc2a9d2a15613d202,
        64'h531bfa5aab4b9a2a,
        64'h09aba94bd15a535a,
        64'haaa3aaa9afaab92b
        },
        {
        64'h8aa92aa8eaa074fe,
        64'ha6d1964514210aad,
        64'ha02aa0ae32b7e280,
        64'hf211b05d2837e402
        },
        {
        64'hc4a86ea9aea6840c,
        64'h92825edaca2a51aa,
        64'h399aabcbaa62802b,
        64'h42af68482a4a3a1a
        },
        {
        64'hb6ea2aa92aabb2be,
        64'ha087a492a552b54b,
        64'h2063a06aaa2ba8ae,
        64'h2d5bf5569053b06a
        },
        {
        64'had6b3d282aa5ee8f,
        64'ha68bb68aa48b24eb,
        64'ha2cab09b268ab28e,
        64'h4aa9eaaaab4b284a
        },
        {
        64'h82ba924aa02d92b1,
        64'ha977992ea93e93b7,
        64'h5052830aabab09a8,
        64'hbaa9aaa860a2f4d7
        },
        {
        64'hb80a2a0129ad73e4,
        64'h73aaf4a2b5aab3e1,
        64'h9b5349456b66a12b,
        64'h6aaf6ea272d7ca52
        },
        {
        64'ha412a154a8285e1c,
        64'ha8422d2aa4aca4ae,
        64'h895524b4b2a51283,
        64'h4aaaaa95a0c1aa45
        },
        {
        64'h9abe0aa9a2ae66aa,
        64'h855bb40a8a3882ab,
        64'h28aaaa2aa92a254f,
        64'h4aafca818d0a8a0a
        },
        {
        64'h0a10caa028ac6ce3,
        64'ha56649526b43c926,
        64'h8168eb6b812a0d2b,
        64'h2aa5d579552b4162
        },
        {
        64'hd4a5950295523a04,
        64'h905792c7b2a3b2aa,
        64'h1d4ad00282029143,
        64'h0aac2aabaaabb15b
        },
        {
        64'hbaadaaa92aa81277,
        64'ha280004119550811,
        64'ha9aba0ae00ab9281,
        64'h5552359fa9a2e9aa
        },
        {
        64'he4ab60a8aead9e98,
        64'ha65a36cae0ca2223,
        64'h2ccaa96aa92b0b2b,
        64'h0aae612b296aee8a
        },
        {
        64'h20a9aaa82aafbcf6,
        64'hb68fb2caa02aa5ab,
        64'h592be88b2846a52c,
        64'h83d81f4a1a6b3a2b
        },
        {
        64'hb5420da82aaf5ea1,
        64'h9253a54aa1b2aa83,
        64'h12439283c28292c2,
        64'heaaa2aab294ba952
        },
        {
        64'h9aabb78969a8a000,
        64'h1b2fadafb8afa6ae,
        64'hcad2ea0aab0a2b2b,
        64'heab62a29ec9128a2
        },
        {
        64'h2a426ad14a8b3bdc,
        64'hccaae886a953aa54,
        64'h584b404b5a2b28ab,
        64'haaa8a5a8c003d242
        },
        {
        64'hb14e2d2028a86af8,
        64'ha92ba16e916fb262,
        64'h049590b682ecab26,
        64'haaa8ea32b4d49594
        },
        {
        64'hd27f52e82aacf295,
        64'h86eba66ab66bd26f,
        64'h32aaa02aa3e3a606,
        64'haaacaaabe3ca922a
        },
        {
        64'h51525261a4ab8086,
        64'haa96ea525b4bd32b,
        64'h112294a682aa4297,
        64'hcaaf9d5ed507555b
        },
        {
        64'hd0a694869557741e,
        64'hd9daa28eaa8abaae,
        64'hb142c24b855b1113,
        64'h2aaaeaaba2aab11a
        },
        {
        64'h82adaaa82aa9b6d6,
        64'ha095364504550ab1,
        64'h282ba0af10af4281,
        64'h7011705fa02be02b
        },
        {
        64'haaaba028aaac54e6,
        64'hd55b5553d44602af,
        64'h00468153d1526553,
        64'h6aa3659ab88b3aab
        },
        {
        64'h20a82aaa2aa590c0,
        64'had1ba2daa36aa12b,
        64'h0a2ba8aa284b294b,
        64'h455b954b2a8a0aaa
        },
        {
        64'ha8a9a0a82aad4aa6,
        64'hd25b866aa12a002b,
        64'haa4facdbb6dbd65a,
        64'h4aaeeaaa2adbaa92
        },
        {
        64'h90a31539a0283e93,
        64'ha9279b2aa92b14a7,
        64'h9952a18aa8aaa80a,
        64'h2aa7eab936924452
        },
        {
        64'hb41a7448cd516dc6,
        64'ha2ab92a2960f943e,
        64'hd446680f2a0baaaa,
        64'h0aae21295543d435
        },
        {
        64'haf17257728a9d2e3,
        64'hafab25aeb594a356,
        64'h2d0535a5a2ada72b,
        64'h8aa9a756ad95aab4
        },
        {
        64'haaa2c000aaadeeba,
        64'hd0569156808382ab,
        64'h280a8553c1931456,
        64'hcaa9caa3aaaa2aaa
        },
        {
        64'h00cad86222abd8ff,
        64'hea57ead252c3d4d3,
        64'h54ab9aab8a4b0a53,
        64'hcaab411dc85a54a2
        },
        {
        64'ha820242a55752e30,
        64'hb46aa26baa2aab2a,
        64'h286ba46ab0cab4cb,
        64'h2aadeaaaaaaaaa2b
        },
        {
        64'ha981aaa9aaa9389a,
        64'h9dedb54931402d09,
        64'h28aaa2afb5a381ed,
        64'hd5746155a857a8aa
        },
        {
        64'h855b65c92aa84888,
        64'h92961253d242554a,
        64'h9497a493a2a32a23,
        64'h0aa96aaab54a3556
        },
        {
        64'h28aaaaa82aa5ccde,
        64'had5bed9aaecba92a,
        64'h0a2be8aaa8ea294b,
        64'he52dedd86c8b8a2b
        },
        {
        64'h95520d0aaaa9bc9a,
        64'h82a2a54aa5238503,
        64'h83578002c283a2aa,
        64'haaaeaaaaad162956
        },
        {
        64'h92a9a7a929ab3a01,
        64'h9baea5aea8aea6ae,
        64'hcad3e24baa4a8b28,
        64'h6a85aa2ae8c12aa2
        },
        {
        64'ha5562551e90befc0,
        64'ha0aba2ae80a29102,
        64'h555751962aa622ae,
        64'h0aa1a8a8b02a5456
        },
        {
        64'haa96aabd2aee9ffb,
        64'h282aa222a807ab62,
        64'h168792ac9208300b,
        64'h4aaba1542418b6b4
        },
        {
        64'h92df8aa1a2a9f6e5,
        64'h957ba6caa6cdd6ca,
        64'h2aaaaaaaaa2b254e,
        64'haaaa082a08bbc28b
        },
        {
        64'h5468d6aa24a4f4b0,
        64'ha90eaaba2a2bd56a,
        64'h700f90a7a0aa212e,
        64'hcaa8d01954065056
        },
        {
        64'hcaae028f551df62a,
        64'h9346935699629baa,
        64'h180a955294538252,
        64'hcaaf6aab2fa998ab
        },
        {
        64'hbaac2aa9caaa31a9,
        64'h84d0944510441825,
        64'he8aba0aa88a39281,
        64'h9813241d20a7e0a3
        },
        {
        64'hfc6828292aa27c98,
        64'h940a5aaa9b2b41ab,
        64'h1ab38a934a53c869,
        64'haaac2a3b2a5a7273
        },
        {
        64'h292baaa82aacae9d,
        64'had1ba4caaccaa96b,
        64'h88abe8cb28cba8ab,
        64'hc13b4d6868ab68aa
        },
        {
        64'h942aba4aaaaa6db0,
        64'h8e8282a6945b956a,
        64'ha48394d684d68653,
        64'haaaf2aaba4aa14a2
        },
        {
        64'h9520a4a9202ca4fc,
        64'h092e9c6aba2b352a,
        64'h0193e8aba92b292a,
        64'h6aabea9a22534317
        },
        {
        64'hb0466a004a917dc1,
        64'haaab88869106917c,
        64'h51624a4b2a2baaaa,
        64'h6aa9a5a85412d554
        },
        {
        64'ha947ab45aae9bfbf,
        64'hab42292eadada895,
        64'h141290a996a8909a,
        64'h4aade2d02a40a30c
        },
        {
        64'h2487b4a8aaa89ab2,
        64'ha8d2a808ac802487,
        64'ha0a8a98aa01bb0c7,
        64'haaa2aaab06aa64aa
        },
        {
        64'h55aa54ab2eae01cc,
        64'hfa47db22d693d60a,
        64'h9090949786f73a57,
        64'heaa8b82920971797
        },
        {
        64'hd557155455561213,
        64'h8403a62ba2a6b782,
        64'h3552e50b8083c863,
        64'h8aaaeaa928aba55a
        },
        {
        64'hbaadaaa86aaa7412,
        64'h8a95874115002295,
        64'haa2aa3aaaaae1284,
        64'hb227f1fc2982632b
        },
        {
        64'hb14b5228aaabdae0,
        64'hc52344129683360a,
        64'h02d3aa53aa4aa92a,
        64'h6aafacab9403b083
        },
        {
        64'ha48a2aa92aaafacd,
        64'hb6b7b6b2a726a482,
        64'h802ba24ba2132756,
        64'ha7f89794929a0a2b
        },
        {
        64'ha6aa88e92aaf76c3,
        64'h92d792178553952a,
        64'h2a4a8a4a8aca92d2,
        64'h2aa02aaaad5b9b4b
        },
        {
        64'hab6b2b0b292fd5ba,
        64'hba4fba7eab6f2b2e,
        64'h053ab9aaa9ab2a8b,
        64'hdaa54a2925a8e02a
        },
        {
        64'h8c8fa201aba199b2,
        64'h692aa1a285ae9dac,
        64'hcb4049554527eb2a,
        64'h0aae6aa33ad28a50
        },
        {
        64'h942eb22368ae92b3,
        64'ha16b256ea96a052a,
        64'h80d682d28a7c292f,
        64'heaad6319214500d6
        },
        {
        64'hb6979689a2ad2481,
        64'hb012ac98a4932696,
        64'h80aa28aaa8233526,
        64'heaada2a900aad0aa
        },
        {
        64'h550a55ab34ab13d2,
        64'hf6d6d69356cad60b,
        64'h92d48896a81704d7,
        64'heaa7894f08571356
        },
        {
        64'hea97c61655d1b40e,
        64'hd113802aa2a2aa93,
        64'ha11bed7bff731063,
        64'h0aab6aaa2aaa2a9b
        },
        {
        64'haa552aa8aaafd9e4,
        64'hb0dcb49914d433d1,
        64'ha8abaa2ba96bb3f9,
        64'h1554e557ad52292b
        },
        {
        64'h952a986a2aacb790,
        64'hca2f5b56c3574916,
        64'hb0ba885a895a4b6a,
        64'haaaeabeb354a3523
        },
        {
        64'ha8a92aabaaa97ec3,
        64'hb4daa64aa36a992b,
        64'h8a2beb6b2f1e2dbb,
        64'h257a1d556a9baa2e
        },
        {
        64'haa0a2b8beaa9765a,
        64'h86a6ae62ac4aa912,
        64'h316a88cb40cf6eee,
        64'haaa86ab9282a812b
        },
        {
        64'h90a215a9a02a3c66,
        64'ha926992aa93f928e,
        64'h5912a9aba92b0909,
        64'h9aa42aa9b283c653
        },
        {
        64'h2845a9436bc6d3c5,
        64'h682aa8aaa88aa8a9,
        64'hd4c750565055c946,
        64'hcaacaaabaaabd207
        },
        {
        64'hb0aa2d5cab2cad88,
        64'ha803250a90ab36ab,
        64'ha9542c34a6ac3caa,
        64'h3aad2aa9aaaca85b
        },
        {
        64'h548bd16bbaa83e92,
        64'hb042b0ca902b54a2,
        64'h2096a196a8d7a057,
        64'h0aaa8ac32a4b8053
        },
        {
        64'h2ab22aab2aaca2b7,
        64'haa53d152d5bad2b3,
        64'h9a1a8942aa222a93,
        64'h0aaf4d2a800a12aa
        },
        {
        64'haa07a9161d53303b,
        64'hd18390a28292aada,
        64'h8d6bad6b80621123,
        64'heaafaaa8aaa9a92a
        },
        {
        64'h2a4c2aa9aaa04ea5,
        64'hb4959415361184a9,
        64'haa2ba22a22aa00a1,
        64'h714022562a9720c2
        },
        {
        64'hf86a682a2aaf12f2,
        64'h812b1962905b448a,
        64'h12b29a92c2d350cb,
        64'hcaa82a9a083a3272
        },
        {
        64'hab4aab29eaa98297,
        64'h9553974a926bdb4a,
        64'h22eb84c2a0c61052,
        64'hd63f905a48ba00ea
        },
        {
        64'h80a8aaca2aabb2ed,
        64'h92860296955a954a,
        64'h896aa94ba0d30296,
        64'h0aacea2a25573643
        },
        {
        64'h21a835a8a12d9902,
        64'h19b6899ead8725af,
        64'hd64bc22baaba88bb,
        64'h3a926aab6a18724f
        },
        {
        64'ha8522c536a4cadbe,
        64'h5caaeeb2ac17281e,
        64'h544b585b5a58da2a,
        64'h2aab2caa76ab52e2
        },
        {
        64'ha8cfaf462928f1ff,
        64'ha123252eb5a7a4e4,
        64'ha4c680c88a64212b,
        64'h2aaf6a552ad424d4
        },
        {
        64'hda3ecb29aaaea4e0,
        64'ha87aae6aa26a826a,
        64'hab25b52295dbe89a,
        64'h6aacaaaaabcb20ab
        },
        {
        64'h0512153ba0ae848e,
        64'hb562d12acabaaaf2,
        64'hdb53890692a682ab,
        64'h2aa9aaabe2aac04a
        },
        {
        64'hd2ab308d15544828,
        64'h929692469a8a12ab,
        64'h844b815384520253,
        64'heaaceaa8aca8022a
        },
        {
        64'haaa8baa96aa54cca,
        64'hb4a5a5cd1404254d,
        64'h2aabaa2f3ea7d684,
        64'h7505a9552a176a4f
        },
        {
        64'h960aa1292eac1bab,
        64'hd12a550e948f16ab,
        64'h12cbaa42aa4a404a,
        64'h6aabaaa9b81630c2
        },
        {
        64'hadabaaa9aaa8a6ce,
        64'hb517b1d69897ccab,
        64'h04aaa52aa9272116,
        64'h865ef40310a380ab
        },
        {
        64'haaa1a06a2aad3ed0,
        64'hd2d2925a954a092a,
        64'h906b888a949386d6,
        64'h0aab6ae8aa038b02
        },
        {
        64'h8a52b1082a2f9dc7,
        64'h3917a93ead379896,
        64'h533ad34bab23892a,
        64'h9aaaaba8f48a1497
        },
        {
        64'h2893a9d42b4a7bfe,
        64'h622aa2aaa28aa929,
        64'hd432555345524142,
        64'h0aa76aab2aabda93
        },
        {
        64'h8552a571a8e8d7e1,
        64'hb646b6949ac62a65,
        64'hb8b5949596143676,
        64'heaa8e4573c543d8d
        },
        {
        64'h92c2f4ab2aac52f1,
        64'hb083acc2a68db696,
        64'ha420a19790b22097,
        64'heaa9282a062b1222
        },
        {
        64'h553ad59bb4ab99b1,
        64'ha2b22ada6a42d10a,
        64'h48a1d0a212af122f,
        64'h0aa5c0595143514b
        },
        {
        64'ha8d4a4540f544249,
        64'h58b392938286aa82,
        64'h8c6bc0739ae318f1,
        64'haaad2aabaaa8a92b
        },
        {
        64'haaacaaa94aa8343e,
        64'ha4851751045582a5,
        64'ha88aa08b30aa1085,
        64'h5406f09f2086e08b
        },
        {
        64'hc16b19c92aaa7cf5,
        64'h9d560b5e992a5102,
        64'h0b2a882ba4ab654a,
        64'h6aacabca9147a942
        },
        {
        64'h26a9aaa8aaa4228e,
        64'hb4b7ba42a32aa58a,
        64'h4aaae81a2a5ba312,
        64'h215cd6140aaa1a2b
        },
        {
        64'hb48922092aafbca7,
        64'hd283902aa1a28522,
        64'h014aa057a2976297,
        64'h6aaaaa28b92a832a
        },
        {
        64'h96abb2ab2aa08fcb,
        64'h1baea1aea4afb6ae,
        64'h6aabeadaaa5b19aa,
        64'haabe6a8b68812aa3
        },
        {
        64'ha958a9526a4359e6,
        64'haaabaeaea4a6ad87,
        64'hc15a4a0b2a8a2a0a,
        64'haaac61aa505b5048
        },
        {
        64'ha956a555aae802e6,
        64'hb6b7b4b4b4b7a916,
        64'h91b495a494b49696,
        64'h8aac351532158091
        },
        {
        64'hd52680ab2aa872e9,
        64'ha8d3a282aa8bb543,
        64'hb426a467a97fad57,
        64'heaac2808f55a34b2
        },
        {
        64'h22ab07682ea31de1,
        64'ha96ad16ac26bcaea,
        64'h2b52a497a6a62026,
        64'hcaa9a8a86aaa2a43
        },
        {
        64'ha02b25ab55713475,
        64'hb0caaa4baa6aa86a,
        64'hd2cb8acab1dab2ca,
        64'h2a8c2aa828a9006b
        },
        {
        64'ha2892aaaaaaa7b8c,
        64'hb4a4b5252d04a5d9,
        64'haa0aa142a51716b5,
        64'h331574142ab228ab
        },
        {
        64'ha18a566baeaf928a,
        64'h8bd227d7a7b63f9a,
        64'h33ebbdebe3eaeb2a,
        64'heaa86daab4ab33aa
        },
        {
        64'hb94aaaabaaaed092,
        64'ha496b6569142914a,
        64'hc0aba123a8aaa88f,
        64'h4559d55010d2101a
        },
        {
        64'hab62aa4a2aaab4a0,
        64'hd29312d2944ab84a,
        64'ha406a6c202921296,
        64'h4aaeaaab2c2aa4a2
        },
        {
        64'h80a986a92aa34848,
        64'h99aea5aeacae36af,
        64'h6a0aea4aaa5b89aa,
        64'h8abbaa8aea432aa2
        },
        {
        64'ha5572551ed411d9b,
        64'h58b3a8d6aa56a917,
        64'h545756d456d5dc97,
        64'h2aaa65aad5aed48f
        },
        {
        64'ha496aa112aaa22e6,
        64'ha56a95299525ab37,
        64'h89b491b5859084ca,
        64'h2aae25203d8ca933
        },
        {
        64'haca63da9aaad70d8,
        64'ha8c2a92ca8aeaca6,
        64'ha0a5a183a0c330dc,
        64'heaa8aaab44aa24ab
        },
        {
        64'h522acaa9a6aa0a02,
        64'haa6ac86a516bd02b,
        64'ha802ac12aca22a0b,
        64'h8aafaae8284e2816
        },
        {
        64'haa02ab440d57f447,
        64'h548294daa2c32a4a,
        64'h8122d92ac3839183,
        64'heaa1eaa8aaaa28ab
        },
        {
        64'hac69baa96aa3399b,
        64'haaa4a8ada505b44d,
        64'h2b2aa92ba8aad680,
        64'hd5576b582b5aeb2a
        },
        {
        64'h845a0f582ea88687,
        64'hd12655b69492745b,
        64'h0242aa52ab2b2b2a,
        64'h6aad2ad9b55b3052
        },
        {
        64'h2b4aaaaaaaa5b79c,
        64'hac17a89aa8832b6a,
        64'hb8aee8cba85e289a,
        64'hc3991da8d82ad8a7
        },
        {
        64'hbaa880192aaa68e3,
        64'h8a138433950214a3,
        64'h244a80d382d30ad6,
        64'h0aafeaa8260b146b
        },
        {
        64'hab4b302b21295348,
        64'h2a9faa6eab5f2a4f,
        64'h152b99aba9aa2a88,
        64'h8ab52aa8b0ab4516
        },
        {
        64'h998a2003caf6d71d,
        64'h2aaaa2a68006817e,
        64'hf15a6a4b2a0aaaaa,
        64'haaa865a9d512d554
        },
        {
        64'ha947aa142aad9296,
        64'haa4f292a29a4aa84,
        64'h98ab90a990a9885a,
        64'h2aab2084b255b805
        },
        {
        64'h8aaae28aaaa81c84,
        64'hd456a052aa81aaaa,
        64'h2aa9a15b957395da,
        64'h6aa862aab2ab22ab
        },
        {
        64'h544ad44a22a935d5,
        64'ha043d4dacadaaada,
        64'hf241a2a282aa824a,
        64'heaa39a2598aab88b
        },
        {
        64'ha8a9a4a915b06e0b,
        64'ha26baa6bab2b292a,
        64'h286aa04ba06bb66b,
        64'hc2a8eaaaaaa8202a
        },
        {
        64'h22813aa96aadcd9d,
        64'hb49512913528a149,
        64'haaaba95ba552d495,
        64'h73537565aaa22aab
        },
        {
        64'hacab82d8aaacdcb3,
        64'he52355069492348b,
        64'h9a42a1528952456a,
        64'h6aa8ae7ab22ab203
        },
        {
        64'ha9aaaaab2aaa98ca,
        64'hb1579152a32ba12a,
        64'h78aba92bac83ac97,
        64'h757a541596ab182a
        },
        {
        64'ha4ab80ab2aaaa29e,
        64'h9a72927294738c0a,
        64'h2ad398d28ab38ae2,
        64'h8aae6aabaad2aadb
        },
        {
        64'h942aa489a1a815b1,
        64'ha22f806ab523152a,
        64'ha113a9aba92aaa2a,
        64'h9aa16a9a22536316
        },
        {
        64'hb6baa26b2aa01ba1,
        64'h286ba122852f35a8,
        64'h69554d450107e36a,
        64'h6aaeeaa34a520b51
        },
        {
        64'ha40b28466a28a430,
        64'ha926b4ae26a8348b,
        64'ha824a8a4acacaa0f,
        64'h8aabea972a54a812
        },
        {
        64'hc95211282baf4dd7,
        64'ha54ea8a2aa90ea52,
        64'hb2699146d5261552,
        64'h4aaf0aa934abb0a3
        },
        {
        64'h49c95b2ba8abc89e,
        64'ha962ed4a6d838d92,
        64'h14c9c2c3ae6aab02,
        64'h8aa8472c474b664a
        },
        {
        64'haa462b470955ea61,
        64'h5592948282872acf,
        64'h41269b0ac203c182,
        64'heaa7eaa82aa928aa
        },
        {
        64'hab992aabaaaaf6a9,
        64'h84a4a50521e5a955,
        64'h3a4b99569096d6b4,
        64'hb1b4a40028b2fa22
        },
        {
        64'ha34ac8aaaeab89b8,
        64'haa5710d6e8c626ff,
        64'ha46aa56be92a6822,
        64'h8aad6f2b152b182a
        },
        {
        64'ha4aa2aaaaaaa9fa5,
        64'had0bad4ab96b91ab,
        64'h0a2a8baa88aaab4e,
        64'hef4fde1c8abb0a4b
        },
        {
        64'ha9522a0baaab1c49,
        64'hcaa20e8abe432903,
        64'h906a9263daf6caa7,
        64'heaa7aaa9a92c012f
        },
        {
        64'h2829ae6aa9291db5,
        64'h1b2e3b2aab2baa2a,
        64'he22af229aa3bba29,
        64'h5abc6a28ecaa282a
        },
        {
        64'h20a7a1516a093be9,
        64'h622aa2aab0aea8a4,
        64'h50b355964453c143,
        64'hea876aaa2aaf4a84
        },
        {
        64'ha8562916aae8e7ae,
        64'h2a432b6ea926a8ac,
        64'h920a92b894a990ab,
        64'h6aab61382088ba4c
        },
        {
        64'ha28252abaaad48b0,
        64'hc157954294a290a2,
        64'ha8a28156a9568817,
        64'h6aa88a802aaaa2ab
        },
        {
        64'h4aabaaa92aa744db,
        64'haa12c862d56ad4aa,
        64'ha893a812a842aa43,
        64'h0aaa62a8ba8eaabb
        },
        {
        64'h9514d555d1597278,
        64'hc662b22fa2a7aad7,
        64'h355ae452d6820603,
        64'haaa7eaabae2ba44a
        },
        {
        64'h2855baa82aabbee8,
        64'ha8a8a8a92555bd51,
        64'ha82aa82b2903b0a8,
        64'hfc416d452a33ea8b
        },
        {
        64'hd4a945abaeaf6c06,
        64'ha92f276ab26b6a6a,
        64'ha88ba0cba80aab29,
        64'h2aabaa6a2a4bea8a
        },
        {
        64'hb24b2aa9aaa7b2dd,
        64'ha496a456a45ba60a,
        64'h6a2ba12aac222484,
        64'ha55ad515030a2a0a
        },
        {
        64'ha308a068a8a9a807,
        64'hdaa34a8a92e38403,
        64'h06d682a69aa70ab6,
        64'h0aaf2aa9216ea87e
        },
        {
        64'h90219118a22ae6b2,
        64'hab36ad6abc0a18b7,
        64'hd543e96bab0a2a2b,
        64'hfaafeba9b08b1532
        },
        {
        64'ha523a521a18d3bcd,
        64'h686ab2aaa96aa14e,
        64'hc9354d614d6fc16b,
        64'haaa92ba0cb53c9ce
        },
        {
        64'ha04eaaacaaab081a,
        64'haa2ab2acb490ab57,
        64'ha4aca8ada948ab4b,
        64'haaa9a856a955a0b4
        },
        {
        64'h9af69e99aaaa5ee6,
        64'hb3d3a0dab2ea9a66,
        64'haa2aaa2aa9031516,
        64'h8aaeeaaa4e130eab
        },
        {
        64'h4a53c2c1aeab6094,
        64'heb56cb43c90acb42,
        64'hd56180aea0af2262,
        64'hcaa5172d550f41a3
        },
        {
        64'hd517155555501621,
        64'h89438006aa87aa97,
        64'h3553c48381a3992a,
        64'h8ab16aaba3aba15a
        },
        {
        64'ha0a1aaaaaaa9b0f0,
        64'hadacb96d2564a121,
        64'h294fb5ae94b704a1,
        64'h7937f8adaa97a856
        },
        {
        64'hb05b4a99aaa9869a,
        64'heb424a56a2562a43,
        64'h00aa80ab8542255b,
        64'heaaa6d6b1d4b2922
        },
        {
        64'ha80b2aa9aaaea4c1,
        64'ha497a4d6bd56a52a,
        64'h28a2e6aa28ab20ae,
        64'h2559155614bba40b
        },
        {
        64'hb40a29a8aaa92a3e,
        64'h9a9a128292a316a3,
        64'ha08ba6b392939282,
        64'h0aa96aabab63aad3
        },
        {
        64'h82aaba992aa91183,
        64'h0d16992ea12b30af,
        64'he8abeb0aab2b094a,
        64'hcaae6aba64522496
        },
        {
        64'hb4ab65506a53cfef,
        64'h422a92aa82aae429,
        64'hb0926ad268535242,
        64'hcaadaaab16a2d494
        },
        {
        64'h968ba4b7a8295c81,
        64'h25aba4a49697b65a,
        64'hac94a424a2042822,
        64'h2aa8235628b4a823
        },
        {
        64'ha2ab00a82aabcca8,
        64'hb157f14a90aa92a2,
        64'ha816a116a4961057,
        64'heaaae8b2288aaaaa
        },
        {
        64'h54c2d8d9b2af1c9a,
        64'ha2d2aac26ad2d04b,
        64'h84a9d2aa1a0b820b,
        64'h2aa3154cb5639007
        },
        {
        64'hc2a95042d5549c38,
        64'hdb5aabcaab2aab2b,
        64'h314bda0acb5b535b,
        64'h4aaa6aaba6a9330b
        },
        {
        64'haa612aa86aa8ac68,
        64'h829524d534a91149,
        64'h22ebb26b2aa302a1,
        64'h55443b452ad322c3
        },
        {
        64'h8b2babe92aaf6893,
        64'h835a515ed3574a2e,
        64'hb81aa34ae962a96b,
        64'h0aa9e9ab8d2a382a
        },
        {
        64'ha94a2b282aab41bb,
        64'h9166b126a923e92a,
        64'h88eb8852845f9542,
        64'h46eafaa982b208ea
        },
        {
        64'h9d430d682aa94886,
        64'hd4428546a8932bcb,
        64'h90568086d2a2528b,
        64'h6aa92aab285f2853
        },
        {
        64'ha8520288232365db,
        64'ha9b6b4cebd0fad5f,
        64'h542af26bab4baa0b,
        64'h8aaf2bab65225587
        },
        {
        64'hb24a26806a818be8,
        64'h6eabbc838d46bb64,
        64'h42d6534a494beaab,
        64'haaadeea8f29256c4
        },
        {
        64'ha8d7aa146aa9cdb1,
        64'haa432b6e292728a6,
        64'h140392a896a81082,
        64'h4aa2637a388c380e
        },
        {
        64'h8aa9f22baaae2a99,
        64'hf15ea544a012ca92,
        64'h392896ea94dad45f,
        64'heaac0aa8baab302b
        },
        {
        64'h4aeaaae822ad6683,
        64'hab6aca6a546bd0eb,
        64'hac0ba9a3aa03a952,
        64'haaa9956bdaff0c3a
        },
        {
        64'hb4a995aa55f6d632,
        64'h9adbaa4aa96ba82a,
        64'hf2db82dabadabada,
        64'h8aa4aaa82029b14b
        },
        {
        64'ha9492aabaaa968d7,
        64'ha949b51134518959,
        64'ha02a96afb4aa05a9,
        64'h38a27a1428562837
        },
        {
        64'h83aa46a8aaab79b9,
        64'h92d25a9eeeb73b73,
        64'h2c4aa96ba92b0a2a,
        64'h0aac25ab392ba86a
        },
        {
        64'haca82aa82aa8adcb,
        64'ha96ab86ab06ab0aa,
        64'h5a2aabaa39ae286e,
        64'he168585e1aba1a0b
        },
        {
        64'h0000000000000000,
        64'h0000000000000000,
        64'h0000000000000000,
        64'h0000000000000000
        },
        {
        64'h0000000000000000,
        64'h0000000000000000,
        64'h0000000000000000,
        64'h0000000000000000
        },
        {
        64'h0000000000000000,
        64'h0000000000000000,
        64'h0000000000000000,
        64'h0000000000000000
        },
        {
        64'h0000000000000000,
        64'h0000000000000000,
        64'h0000000000000000,
        64'h0000000000000000
        },
        {
        64'h0000000000000000,
        64'h0000000000000000,
        64'h0000000000000000,
        64'h0000000000000000
        },
        {
        64'h0000000000000000,
        64'h0000000000000000,
        64'h0000000000000000,
        64'h0000000000000000
        }
    }
    // dont open if you dont know what it means
)
(
    input clk,
    input rst,
    input [$clog2(NUM_AXONS)-1:0] axon_number,
    input [$clog2(NUM_NEURONS)-1:0] neuron_number,

    output matrix_connection
);
    
    // wire output_matrix_connection;
    wire [NUM_NEURONS-1:0] neuron_con_outs;

    // instance of 256 neuron connection
	genvar curr_neuron_num;
	
	for (curr_neuron_num = 0; curr_neuron_num < NUM_NEURONS; curr_neuron_num = curr_neuron_num + 1) begin 
		neuron_con #(
            .NUM_AXONS(NUM_AXONS),
            .LUT_INIT(LUT_INIT[curr_neuron_num])
        ) neuron_con_inst (
            .clk(clk),
            .rst(rst),
            .axon_number(axon_number), 
            .connection(neuron_con_outs[curr_neuron_num])
        );
	end


    // // mux logic
    // always @(posedge clk) begin
    //     if (rst)
    //         matrix_connection <= 1'b0;
    //     else begin
    //         matrix_connection = neuron_con_outs[neuron_number];
    //     end
    // end

    assign matrix_connection = neuron_con_outs[neuron_number];
endmodule